module trade_SMA #(
    // makes it adjustable from TLU
    parameter data_width = 16,
    parameter [data_width:0] threshold = 17'd4928,  
    parameter [1:0] confluence_threshold = 2'd3
)(
    input logic clk,
    input logic rst,
    input logic data_valid_pre,
    input logic[data_width-1:0] data_5,
    input logic[data_width-1:0] data_10,
    input logic[data_width-1:0] data_20,
    input logic[data_width-1:0] data_50,
    input logic[data_width-1:0] data_100,
    input logic[data_width-1:0] data_200,
    output logic buy_signal,
    output logic sell_signal,
    output logic data_valid_sma
);


    logic [data_width-1:0] prev_5, prev_10, prev_20, prev_50, prev_100, prev_200;
    logic rising_5, rising_10, rising_20, rising_50, rising_100, rising_200;
    logic falling_5, falling_10, falling_20, falling_50, falling_100, falling_200;
    logic [data_width:0] up_score, down_score;
    
    logic strong_uptrend, strong_downtrend;
    logic confluence_rising, confluence_falling;

    logic buy_signal_next, sell_signal_next;

    // getting previous SMA values for trend detection
    // can be made to look more clean with registers if needed
    // but FPGA compiler should be able to optimise this

    always_ff @( posedge clk ) begin
        if (rst) begin
            prev_5 <= {data_width{1'b0}};
            prev_10 <= {data_width{1'b0}};
            prev_20 <= {data_width{1'b0}};
            prev_50 <= {data_width{1'b0}};
            prev_100 <= {data_width{1'b0}};
            prev_200 <= {data_width{1'b0}};
        end
        else begin 
            prev_5 <= data_5;
            prev_10 <= data_10;
            prev_20 <= data_20;
            prev_50 <= data_50;
            prev_100 <= data_100;
            prev_200 <= data_200;
        end  
    end 

    always_comb begin
        rising_5   = data_5   > prev_5;
        rising_10  = data_10  > prev_10;
        rising_20  = data_20  > prev_20;
        rising_50  = data_50  > prev_50;
        rising_100 = data_100 > prev_100;
        rising_200 = data_200 > prev_200; 

        falling_5   = data_5   < prev_5; 
        falling_10  = data_10  < prev_10;
        falling_20  = data_20  < prev_20;
        falling_50  = data_50  < prev_50;
        falling_100 = data_100 < prev_100;
        falling_200 = data_200 < prev_200;        
       
    end

    //implementing scoring system for trend strength
    assign up_score   = (data_5 - data_20) + (data_10 - data_50);
    assign down_score = (data_20 - data_5) + (data_50 - data_10);
    assign strong_uptrend   = up_score > threshold;
    assign strong_downtrend = down_score > threshold;


    // confluence detection
    always_ff @( posedge clk ) begin 
        if (rst) begin
            confluence_rising <= 1'b0;
            confluence_falling <= 1'b0;
        end
        else begin
            // counting how many SMAs are rising/falling
            confluence_rising <= (rising_5 + rising_10 + rising_20 + rising_50 + rising_100 + rising_200) >= confluence_threshold;
            confluence_falling <= (falling_5 + falling_10 + falling_20 + falling_50 + falling_100 + falling_200) >= confluence_threshold;
        end
    end

    // generating buy/sell signals based on trend strength and confluence
    assign buy_signal_next  = strong_uptrend && confluence_rising;
    assign sell_signal_next = strong_downtrend && confluence_falling;
    

    // synchronising the signals for TPU
    always_ff @( posedge clk ) begin 
        if (rst) begin
            buy_signal  <= 1'b0;
            sell_signal <= 1'b0;
        end
        else begin
            buy_signal  <= buy_signal_next;
            sell_signal <= sell_signal_next;
            data_valid_sma <= data_valid_pre;
        end
    end
    

    

    
endmodule

