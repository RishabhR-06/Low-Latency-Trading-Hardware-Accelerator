module sqr_root #(
    parameter[5:0] size = 5'd16,
) (
    input logic clk,
    input logic rst,
    input logic[size-1:0] data_in,
    output logic[size-1:0] rooted_data_out
);


    //square roots the input data
    //researching algorithims for now



    
endmodule